library verilog;
use verilog.vl_types.all;
entity folder_tb is
end folder_tb;
